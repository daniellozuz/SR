module adder_latency0
(
	// input ports
	input [7:0] a,
	input [7:0] b,
	// output ports
	output [7:0] y
)
assign y = a + b;

endmodule;
