module simple_module
(
	// input ports
	input a,
	input b,
	input [3:0] x,
	// output ports
	output c,
	output [3:0] y
);
// module content
endmodule